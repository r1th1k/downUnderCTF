BZh91AY&SY�5�P �߀Py���߰����P�r":-� 0&&�	�&L�&	����T��@ �  �� SD����I�4ф   4 9�14L�2da0M4����$I�&&F�Sa&ИS�~��4=L�ޤ�n�K!����䯟�Y?�0T*T�U'��%��j��ED�I�$�X�����b�|��4xH�*֡SA=���0��܈"�{�ݜ�M�
t�8�סc��\��4b�ъ�_�4�k ���$�3:LW����4�1�WϩهXk������������n����%�����%NW\-;Z�$��E�"FuR&�9}��\�zO;d˘���!&YRI$�C�����!
�A��3J$�w3`x�A+f�Ƀ�]��W��ֲҙ�iS�R2���Ye3ai������ΣM6�6�叹�\4���f�'絡����~^K�jϜ��]mF�3�P��J+����� , ���E!K����ͩ��=Y���Δש�#���|a�~���Vl����5�{��~���NsІ����G�pT}X>\�ų�8�Y1�R��^-��-DD�Dud�>�������@�B(�����4$�@���f(2$[�5�|�����^���_\��nv[��T���Z{����N-���IeS�y��W��w�/�â(��I��kJ��x�Csw�>�_����5%��(�����v���|�iZ�4��v���}E����d����=�'��9�y�#x�S��,��G*�7�ͧ��l�U����xw���UZ(��;{0��c�w��c��x�IY��MT��J��-݌K��7�y,��V|���Զ�w�`��s��Ҽx�IM3h�����>��d����t���zX�r9����פ<%U�;z�ͥ#����nY�<�S��ɥ�6�:"k�2�F,�uｽ�^���T��NޭF2��;���.y��y���f���w��6���xp\h�P�I�i���ӵi7��wm��Z8��yY?]*�}&��a���ĥ:�'b��W4L����)�ᮢ�